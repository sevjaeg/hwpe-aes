/*
 * mac_engine.sv
 * Francesco Conti <fconti@iis.ee.ethz.ch>
 *
 * Copyright (C) 2018 ETH Zurich, University of Bologna
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 */

import mac_package::*;

module mac_engine
(
  // global signals
  input  logic                   clk_i,
  input  logic                   rst_ni,
  // input a stream
  hwpe_stream_intf_stream.sink   a_i,
  // input b stream
  hwpe_stream_intf_stream.sink   b_i,
  // output d stream
  hwpe_stream_intf_stream.source d_o,
  // control channel
  input  ctrl_engine_t           ctrl_i,
  output flags_engine_t          flags_o
);

  logic unsigned [$clog2(MAC_CNT_LEN):0] cnt;
  logic unsigned [$clog2(MAC_CNT_LEN):0] r_cnt;
  logic signed [127:0] r_word;
  logic signed [127:0] r_key;
  logic signed [127:0] aes_out;
  logic signed [127:0] r_aes;
  logic               r_word_valid;
  logic               r_word_ready;
  logic               r_key_valid;
  logic               r_key_ready;
  logic               r_aes_valid;
  logic               r_aes_ready;
  logic               aes_valid;
  logic               aes_ready;
  logic               aes_start;
  logic               aes_busy;

  aes_cipher_top i_aes(
    .clk (clk_i),
    .rst (rst_ni),
    .ld  (aes_start),
    .done(aes_valid),
    .key (r_key),
    .text_in (r_word),
    .text_out (aes_out)
  );

  // register value updates
  always_ff @(posedge clk_i or negedge rst_ni)
  begin : mult_pipe_data
    if(~rst_ni) begin
      r_word <= '0;
      r_key  <= '0;
      r_aes  <= '0;
    end
    else if (ctrl_i.clear) begin
      r_word <= '0;
      r_key  <= '0;
      r_aes  <= '0;
    end
    else if (ctrl_i.enable) begin
      // updates at valid handshake at input
      if (a_i.valid & a_i.ready) begin
        r_word <= $signed(a_i.data);
      end
      if (b_i.valid & b_i.ready) begin
        r_key <= $signed(b_i.data);
      end
      if (aes_valid & aes_ready) begin
        r_aes <= aes_out;
      end
    end
  end

  // r_word is valid following a valid handshake
  always_ff @(posedge clk_i or negedge rst_ni)
  begin : r_word_val
    if(~rst_ni) begin
      r_word_valid <= '0;
    end
    else if (ctrl_i.clear) begin
      r_word_valid <= '0;
    end
    else if (ctrl_i.enable) begin
      // r_word_valid is re-evaluated after a valid handshake or in transition to 1
      if ((a_i.valid) | (r_word_valid & r_word_ready)) begin
        r_word_valid <= a_i.valid;
      end
    end
  end

  // r_key is valid following a valid handshake
  always_ff @(posedge clk_i or negedge rst_ni)
  begin : r_key_val
    if(~rst_ni) begin
      r_key_valid <= '0;
    end
    else if (ctrl_i.clear) begin
      r_key_valid <= '0;
    end
    else if (ctrl_i.enable) begin
      // r_word_valid is re-evaluated after a valid handshake or in transition to 1
      if ((b_i.valid) | (r_key_valid & r_key_ready)) begin
        r_key_valid <= b_i.valid;
      end
    end
  end

  assign aes_start = r_word_valid & r_key_valid & (~aes_busy);

  // r_aes is valid following a valid handshake
  always_ff @(posedge clk_i or negedge rst_ni)
  begin : proc_aes_busy
    if(~rst_ni) begin
      aes_busy <= '0;
    end
    else if (ctrl_i.clear) begin
      aes_busy <= '0;
    end
    else if (ctrl_i.enable) begin
      // r_word_valid is re-evaluated after a valid handshake or in transition to 1
      if (aes_start) begin
        aes_busy <= '1;
      end
      if (aes_valid) begin
        aes_busy <= '0;
      end
    end
  end

  // r_aes is valid following a valid handshake
  always_ff @(posedge clk_i or negedge rst_ni)
  begin : r_aes_val
    if(~rst_ni) begin
      r_aes_valid <= '0;
    end
    else if (ctrl_i.clear) begin
      r_aes_valid <= '0;
    end
    else if (ctrl_i.enable) begin
      // r_word_valid is re-evaluated after a valid handshake or in transition to 1
      if ((aes_valid) | (r_aes_valid & r_aes_ready)) begin
        r_aes_valid <= aes_valid;
      end
    end
  end

  always_comb
  begin
    d_o.data  = r_aes[31:0];//32'hffffffff; //$signed(r_word);
    d_o.valid = ctrl_i.enable & aes_valid;//r_word_valid;
    d_o.strb  = '1; // for now, strb is always '1
  end

  // The control counter is implemented directly inside this module; as the control is
  // minimal, it was not deemed convenient to move it to another submodule. For bigger
  // FSMs that is typically the most advantageous choice.

  always_comb
  begin
    cnt = r_cnt + 1;
  end

  always_ff @(posedge clk_i or negedge rst_ni)
  begin
    if(~rst_ni) begin
      r_cnt <= '0;
    end
    else if(ctrl_i.clear) begin
      r_cnt <= '0;
    end
    else if(ctrl_i.enable) begin
      if ((ctrl_i.start == 1'b1) || ((r_cnt > 0) && (r_cnt < ctrl_i.len) && (r_word_valid & r_word_ready == 1'b1))) begin
        r_cnt <= cnt;
      end
    end
  end

  assign flags_o.cnt = r_cnt;
  assign flags_o.acc_valid = r_aes_valid;

  // Ready signals have to be propagated backwards through pipeline stages (combinationally).
  // To avoid deadlocks, the following rules have to be followed:
  //  1) transition of ready CAN depend on the current state of valid
  //  2) transition of valid CANNOT depend on the current state of ready
  //  3) transition 1->0 of valid MUST depend on (previous) ready (i.e., once the valid goes
  //     to 1 it cannot go back to 0 until there is a valid handshake)
  // In the following:
  // R_valid & R_ready denominate the handshake at the *output* (Q port) of pipe register R

  assign a_i.ready = (r_word_ready & a_i.valid & b_i.valid) | (~a_i.valid & ~b_i.valid);
  assign b_i.ready = (r_key_ready & a_i.valid  & b_i.valid) | (~a_i.valid & ~b_i.valid);

  // aes accepts if output register free and AES core not busy
  assign r_word_ready = (aes_ready & (~aes_busy | ~aes_start));
  assign r_key_ready = (aes_ready & (~aes_busy | ~aes_start));

  // aes reg accepts if output ready or nothing useful in register
  assign aes_ready =  r_aes_ready | (~r_aes_valid);

  assign r_aes_ready = d_o.ready;
  
endmodule // mac_engine
